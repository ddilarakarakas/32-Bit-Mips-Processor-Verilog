module bus(out,ins,pc);
	output[31:0] out;
	input[25:0] ins;
	input[3:0] pc;
	or(out[31],pc[3],0);
	or(out[30],pc[2],0);
	or(out[29],pc[1],0);
	or(out[28],pc[0],0);
	or(out[27],ins[25],0);
	or(out[26],ins[24],0);
	or(out[25],ins[23],0);
	or(out[24],ins[22],0);
	or(out[23],ins[21],0);
	or(out[22],ins[20],0);
	or(out[21],ins[19],0);
	or(out[20],ins[18],0);
	or(out[19],ins[17],0);
	or(out[18],ins[16],0);
	or(out[17],ins[15],0);
	or(out[16],ins[14],0);
	or(out[15],ins[13],0);
	or(out[14],ins[12],0);
	or(out[13],ins[11],0);
	or(out[12],ins[10],0);
	or(out[11],ins[9],0);
	or(out[10],ins[8],0);
	or(out[9],ins[7],0);
	or(out[8],ins[6],0);
	or(out[7],ins[5],0);
	or(out[6],ins[4],0);
	or(out[5],ins[3],0);
	or(out[4],ins[2],0);
	or(out[3],ins[1],0);
	or(out[2],ins[0],0);
	or(out[1],0,0);
	or(out[0],0,0);
endmodule 